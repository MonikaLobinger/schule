h1, h2, h3, h4, h5, h6 {
  margin-bottom: 0rem;
  margin-top: 0rem;
  padding-top: 0rem;
  padding-top: 0rem;
  margin-block-end: 0rem;
  margin-block-start: 0rem;
}
h1 {
   font-size: 2rem ;
   margin-bottom: 0.5rem;
 }
h2 {
   font-size: 1.5rem ;
   margin-bottom: 0.5rem;
 }
h3{
   font-size: 1.3rem ;
}
p  {
  line-height: 1.3rem;
  margin-top: 0rem;
  margin-bottom: 0.3rem;
}
li {
  line-height: 1.2rem;
}
.el-h3, .el-ul {
  margin: 0;
  padding: 0;
}
