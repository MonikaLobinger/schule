/* Damit das Plugin "Webpage HTML Export" den Dateinamen nicht als H1 anzeigt */
.page-title, .mod-header {
  background-color: red !important;
  display:none;
}
/* Ich verwende viele Links, sie müssen dunkler sein */
body {
    --link-color: #4169E1; /* Internal link color (e.g., royal blue) */
    --link-color-hover: #0000CD; /* Internal link hover color (e.g., medium blue) */
    --link-external-color: #4169E1; /* External link color (e.g., royal blue) */
    --link-external-color-hover: #0000CD; /* External link hover color (e.g., medium blue) */
    --link-decoration: none;
    --link-decoration-hover: none;
}
